// TestRO.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module TestRO (
		input  wire        clk_clk,               //          clk.clk
		output wire [31:0] dacctrl_export,        //      dacctrl.export
		output wire        ext_rst_export,        //      ext_rst.export
		output wire        exttrg_0_export,       //     exttrg_0.export
		input  wire [31:0] fifo_0_in_writedata,   //    fifo_0_in.writedata
		input  wire        fifo_0_in_write,       //             .write
		output wire        fifo_0_in_waitrequest, //             .waitrequest
		input  wire [31:0] fifo_1_in_writedata,   //    fifo_1_in.writedata
		input  wire        fifo_1_in_write,       //             .write
		output wire        fifo_1_in_waitrequest, //             .waitrequest
		input  wire        reset_reset_n,         //        reset.reset_n
		input  wire [31:0] version_info_export,   // version_info.export
		output wire        write_en_export        //     write_en.export
	);

	wire   [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire          nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire          nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire   [29:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire    [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire          nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire          nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire   [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire   [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire          nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire   [28:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire          nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire   [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire   [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire   [31:0] mm_interconnect_0_fifo_0_out_readdata;                       // fifo_0:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_0_out_readdata
	wire          mm_interconnect_0_fifo_0_out_waitrequest;                    // fifo_0:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_0_out_waitrequest
	wire          mm_interconnect_0_fifo_0_out_read;                           // mm_interconnect_0:fifo_0_out_read -> fifo_0:avalonmm_read_slave_read
	wire   [31:0] mm_interconnect_0_fifo_1_out_readdata;                       // fifo_1:avalonmm_read_slave_readdata -> mm_interconnect_0:fifo_1_out_readdata
	wire          mm_interconnect_0_fifo_1_out_waitrequest;                    // fifo_1:avalonmm_read_slave_waitrequest -> mm_interconnect_0:fifo_1_out_waitrequest
	wire          mm_interconnect_0_fifo_1_out_read;                           // mm_interconnect_0:fifo_1_out_read -> fifo_1:avalonmm_read_slave_read
	wire   [31:0] mm_interconnect_0_fifo_0_out_csr_readdata;                   // fifo_0:rdclk_control_slave_readdata -> mm_interconnect_0:fifo_0_out_csr_readdata
	wire    [2:0] mm_interconnect_0_fifo_0_out_csr_address;                    // mm_interconnect_0:fifo_0_out_csr_address -> fifo_0:rdclk_control_slave_address
	wire          mm_interconnect_0_fifo_0_out_csr_read;                       // mm_interconnect_0:fifo_0_out_csr_read -> fifo_0:rdclk_control_slave_read
	wire          mm_interconnect_0_fifo_0_out_csr_write;                      // mm_interconnect_0:fifo_0_out_csr_write -> fifo_0:rdclk_control_slave_write
	wire   [31:0] mm_interconnect_0_fifo_0_out_csr_writedata;                  // mm_interconnect_0:fifo_0_out_csr_writedata -> fifo_0:rdclk_control_slave_writedata
	wire   [31:0] mm_interconnect_0_fifo_1_out_csr_readdata;                   // fifo_1:rdclk_control_slave_readdata -> mm_interconnect_0:fifo_1_out_csr_readdata
	wire    [2:0] mm_interconnect_0_fifo_1_out_csr_address;                    // mm_interconnect_0:fifo_1_out_csr_address -> fifo_1:rdclk_control_slave_address
	wire          mm_interconnect_0_fifo_1_out_csr_read;                       // mm_interconnect_0:fifo_1_out_csr_read -> fifo_1:rdclk_control_slave_read
	wire          mm_interconnect_0_fifo_1_out_csr_write;                      // mm_interconnect_0:fifo_1_out_csr_write -> fifo_1:rdclk_control_slave_write
	wire   [31:0] mm_interconnect_0_fifo_1_out_csr_writedata;                  // mm_interconnect_0:fifo_1_out_csr_writedata -> fifo_1:rdclk_control_slave_writedata
	wire          mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [127:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [14:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [15:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire          mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [127:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire          mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire          mm_interconnect_0_write_en_pio_s1_chipselect;                // mm_interconnect_0:write_en_pio_s1_chipselect -> write_en_pio:chipselect
	wire   [31:0] mm_interconnect_0_write_en_pio_s1_readdata;                  // write_en_pio:readdata -> mm_interconnect_0:write_en_pio_s1_readdata
	wire    [1:0] mm_interconnect_0_write_en_pio_s1_address;                   // mm_interconnect_0:write_en_pio_s1_address -> write_en_pio:address
	wire          mm_interconnect_0_write_en_pio_s1_write;                     // mm_interconnect_0:write_en_pio_s1_write -> write_en_pio:write_n
	wire   [31:0] mm_interconnect_0_write_en_pio_s1_writedata;                 // mm_interconnect_0:write_en_pio_s1_writedata -> write_en_pio:writedata
	wire          mm_interconnect_0_exttrg_0_s1_chipselect;                    // mm_interconnect_0:exttrg_0_s1_chipselect -> exttrg_0:chipselect
	wire   [31:0] mm_interconnect_0_exttrg_0_s1_readdata;                      // exttrg_0:readdata -> mm_interconnect_0:exttrg_0_s1_readdata
	wire    [1:0] mm_interconnect_0_exttrg_0_s1_address;                       // mm_interconnect_0:exttrg_0_s1_address -> exttrg_0:address
	wire          mm_interconnect_0_exttrg_0_s1_write;                         // mm_interconnect_0:exttrg_0_s1_write -> exttrg_0:write_n
	wire   [31:0] mm_interconnect_0_exttrg_0_s1_writedata;                     // mm_interconnect_0:exttrg_0_s1_writedata -> exttrg_0:writedata
	wire          mm_interconnect_0_dacctrl_s1_chipselect;                     // mm_interconnect_0:dacctrl_s1_chipselect -> dacctrl:chipselect
	wire   [31:0] mm_interconnect_0_dacctrl_s1_readdata;                       // dacctrl:readdata -> mm_interconnect_0:dacctrl_s1_readdata
	wire    [1:0] mm_interconnect_0_dacctrl_s1_address;                        // mm_interconnect_0:dacctrl_s1_address -> dacctrl:address
	wire          mm_interconnect_0_dacctrl_s1_write;                          // mm_interconnect_0:dacctrl_s1_write -> dacctrl:write_n
	wire   [31:0] mm_interconnect_0_dacctrl_s1_writedata;                      // mm_interconnect_0:dacctrl_s1_writedata -> dacctrl:writedata
	wire   [31:0] mm_interconnect_0_version_info_s1_readdata;                  // version_info:readdata -> mm_interconnect_0:version_info_s1_readdata
	wire    [1:0] mm_interconnect_0_version_info_s1_address;                   // mm_interconnect_0:version_info_s1_address -> version_info:address
	wire          mm_interconnect_0_ext_rst_s1_chipselect;                     // mm_interconnect_0:ext_rst_s1_chipselect -> ext_rst:chipselect
	wire   [31:0] mm_interconnect_0_ext_rst_s1_readdata;                       // ext_rst:readdata -> mm_interconnect_0:ext_rst_s1_readdata
	wire    [1:0] mm_interconnect_0_ext_rst_s1_address;                        // mm_interconnect_0:ext_rst_s1_address -> ext_rst:address
	wire          mm_interconnect_0_ext_rst_s1_write;                          // mm_interconnect_0:ext_rst_s1_write -> ext_rst:write_n
	wire   [31:0] mm_interconnect_0_ext_rst_s1_writedata;                      // mm_interconnect_0:ext_rst_s1_writedata -> ext_rst:writedata
	wire          irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire   [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire          rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [dacctrl:reset_n, ext_rst:reset_n, exttrg_0:reset_n, fifo_0:rdreset_n, fifo_0:wrreset_n, fifo_1:rdreset_n, fifo_1:wrreset_n, irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator:in_reset, version_info:reset_n, write_en_pio:reset_n]
	wire          rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset]
	wire          rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [onchip_memory2_0:reset_req, rst_translator_001:reset_req_in]
	wire          nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> rst_controller_001:reset_in1

	TestRO_dacctrl dacctrl (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_dacctrl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_dacctrl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_dacctrl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_dacctrl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_dacctrl_s1_readdata),   //                    .readdata
		.out_port   (dacctrl_export)                           // external_connection.export
	);

	TestRO_ext_rst ext_rst (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_ext_rst_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ext_rst_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ext_rst_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ext_rst_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ext_rst_s1_readdata),   //                    .readdata
		.out_port   (ext_rst_export)                           // external_connection.export
	);

	TestRO_ext_rst exttrg_0 (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_exttrg_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_exttrg_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_exttrg_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_exttrg_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_exttrg_0_s1_readdata),   //                    .readdata
		.out_port   (exttrg_0_export)                           // external_connection.export
	);

	TestRO_fifo_0 fifo_0 (
		.wrclock                          (clk_clk),                                    //    clk_in.clk
		.wrreset_n                        (~rst_controller_reset_out_reset),            //  reset_in.reset_n
		.rdclock                          (clk_clk),                                    //   clk_out.clk
		.rdreset_n                        (~rst_controller_reset_out_reset),            // reset_out.reset_n
		.avalonmm_write_slave_writedata   (fifo_0_in_writedata),                        //        in.writedata
		.avalonmm_write_slave_write       (fifo_0_in_write),                            //          .write
		.avalonmm_write_slave_waitrequest (fifo_0_in_waitrequest),                      //          .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_0_out_readdata),      //       out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_0_out_read),          //          .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_0_out_waitrequest),   //          .waitrequest
		.rdclk_control_slave_address      (mm_interconnect_0_fifo_0_out_csr_address),   //   out_csr.address
		.rdclk_control_slave_read         (mm_interconnect_0_fifo_0_out_csr_read),      //          .read
		.rdclk_control_slave_writedata    (mm_interconnect_0_fifo_0_out_csr_writedata), //          .writedata
		.rdclk_control_slave_write        (mm_interconnect_0_fifo_0_out_csr_write),     //          .write
		.rdclk_control_slave_readdata     (mm_interconnect_0_fifo_0_out_csr_readdata)   //          .readdata
	);

	TestRO_fifo_0 fifo_1 (
		.wrclock                          (clk_clk),                                    //    clk_in.clk
		.wrreset_n                        (~rst_controller_reset_out_reset),            //  reset_in.reset_n
		.rdclock                          (clk_clk),                                    //   clk_out.clk
		.rdreset_n                        (~rst_controller_reset_out_reset),            // reset_out.reset_n
		.avalonmm_write_slave_writedata   (fifo_1_in_writedata),                        //        in.writedata
		.avalonmm_write_slave_write       (fifo_1_in_write),                            //          .write
		.avalonmm_write_slave_waitrequest (fifo_1_in_waitrequest),                      //          .waitrequest
		.avalonmm_read_slave_readdata     (mm_interconnect_0_fifo_1_out_readdata),      //       out.readdata
		.avalonmm_read_slave_read         (mm_interconnect_0_fifo_1_out_read),          //          .read
		.avalonmm_read_slave_waitrequest  (mm_interconnect_0_fifo_1_out_waitrequest),   //          .waitrequest
		.rdclk_control_slave_address      (mm_interconnect_0_fifo_1_out_csr_address),   //   out_csr.address
		.rdclk_control_slave_read         (mm_interconnect_0_fifo_1_out_csr_read),      //          .read
		.rdclk_control_slave_writedata    (mm_interconnect_0_fifo_1_out_csr_writedata), //          .writedata
		.rdclk_control_slave_write        (mm_interconnect_0_fifo_1_out_csr_write),     //          .write
		.rdclk_control_slave_readdata     (mm_interconnect_0_fifo_1_out_csr_readdata)   //          .readdata
	);

	TestRO_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	TestRO_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	TestRO_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	TestRO_version_info version_info (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_version_info_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_version_info_s1_readdata), //                    .readdata
		.in_port  (version_info_export)                         // external_connection.export
	);

	TestRO_ext_rst write_en_pio (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_write_en_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_write_en_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_write_en_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_write_en_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_write_en_pio_s1_readdata),   //                    .readdata
		.out_port   (write_en_export)                               // external_connection.export
	);

	TestRO_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset  (rst_controller_001_reset_out_reset),                          //  jtag_uart_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.dacctrl_s1_address                             (mm_interconnect_0_dacctrl_s1_address),                        //                               dacctrl_s1.address
		.dacctrl_s1_write                               (mm_interconnect_0_dacctrl_s1_write),                          //                                         .write
		.dacctrl_s1_readdata                            (mm_interconnect_0_dacctrl_s1_readdata),                       //                                         .readdata
		.dacctrl_s1_writedata                           (mm_interconnect_0_dacctrl_s1_writedata),                      //                                         .writedata
		.dacctrl_s1_chipselect                          (mm_interconnect_0_dacctrl_s1_chipselect),                     //                                         .chipselect
		.ext_rst_s1_address                             (mm_interconnect_0_ext_rst_s1_address),                        //                               ext_rst_s1.address
		.ext_rst_s1_write                               (mm_interconnect_0_ext_rst_s1_write),                          //                                         .write
		.ext_rst_s1_readdata                            (mm_interconnect_0_ext_rst_s1_readdata),                       //                                         .readdata
		.ext_rst_s1_writedata                           (mm_interconnect_0_ext_rst_s1_writedata),                      //                                         .writedata
		.ext_rst_s1_chipselect                          (mm_interconnect_0_ext_rst_s1_chipselect),                     //                                         .chipselect
		.exttrg_0_s1_address                            (mm_interconnect_0_exttrg_0_s1_address),                       //                              exttrg_0_s1.address
		.exttrg_0_s1_write                              (mm_interconnect_0_exttrg_0_s1_write),                         //                                         .write
		.exttrg_0_s1_readdata                           (mm_interconnect_0_exttrg_0_s1_readdata),                      //                                         .readdata
		.exttrg_0_s1_writedata                          (mm_interconnect_0_exttrg_0_s1_writedata),                     //                                         .writedata
		.exttrg_0_s1_chipselect                         (mm_interconnect_0_exttrg_0_s1_chipselect),                    //                                         .chipselect
		.fifo_0_out_read                                (mm_interconnect_0_fifo_0_out_read),                           //                               fifo_0_out.read
		.fifo_0_out_readdata                            (mm_interconnect_0_fifo_0_out_readdata),                       //                                         .readdata
		.fifo_0_out_waitrequest                         (mm_interconnect_0_fifo_0_out_waitrequest),                    //                                         .waitrequest
		.fifo_0_out_csr_address                         (mm_interconnect_0_fifo_0_out_csr_address),                    //                           fifo_0_out_csr.address
		.fifo_0_out_csr_write                           (mm_interconnect_0_fifo_0_out_csr_write),                      //                                         .write
		.fifo_0_out_csr_read                            (mm_interconnect_0_fifo_0_out_csr_read),                       //                                         .read
		.fifo_0_out_csr_readdata                        (mm_interconnect_0_fifo_0_out_csr_readdata),                   //                                         .readdata
		.fifo_0_out_csr_writedata                       (mm_interconnect_0_fifo_0_out_csr_writedata),                  //                                         .writedata
		.fifo_1_out_read                                (mm_interconnect_0_fifo_1_out_read),                           //                               fifo_1_out.read
		.fifo_1_out_readdata                            (mm_interconnect_0_fifo_1_out_readdata),                       //                                         .readdata
		.fifo_1_out_waitrequest                         (mm_interconnect_0_fifo_1_out_waitrequest),                    //                                         .waitrequest
		.fifo_1_out_csr_address                         (mm_interconnect_0_fifo_1_out_csr_address),                    //                           fifo_1_out_csr.address
		.fifo_1_out_csr_write                           (mm_interconnect_0_fifo_1_out_csr_write),                      //                                         .write
		.fifo_1_out_csr_read                            (mm_interconnect_0_fifo_1_out_csr_read),                       //                                         .read
		.fifo_1_out_csr_readdata                        (mm_interconnect_0_fifo_1_out_csr_readdata),                   //                                         .readdata
		.fifo_1_out_csr_writedata                       (mm_interconnect_0_fifo_1_out_csr_writedata),                  //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),               //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                         .clken
		.version_info_s1_address                        (mm_interconnect_0_version_info_s1_address),                   //                          version_info_s1.address
		.version_info_s1_readdata                       (mm_interconnect_0_version_info_s1_readdata),                  //                                         .readdata
		.write_en_pio_s1_address                        (mm_interconnect_0_write_en_pio_s1_address),                   //                          write_en_pio_s1.address
		.write_en_pio_s1_write                          (mm_interconnect_0_write_en_pio_s1_write),                     //                                         .write
		.write_en_pio_s1_readdata                       (mm_interconnect_0_write_en_pio_s1_readdata),                  //                                         .readdata
		.write_en_pio_s1_writedata                      (mm_interconnect_0_write_en_pio_s1_writedata),                 //                                         .writedata
		.write_en_pio_s1_chipselect                     (mm_interconnect_0_write_en_pio_s1_chipselect)                 //                                         .chipselect
	);

	TestRO_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
