
module ADCINCLKCTRL (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
