
module SYS_GCLK (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
